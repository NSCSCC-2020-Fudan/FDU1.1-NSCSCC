module issue 
    import common::*;
    import queue_pkg::*(
    
);
    issue_queue_t issue_queue; 
endmodule