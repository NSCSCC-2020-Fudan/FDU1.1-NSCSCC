`ifndef DISABLE_DEFAULT_TU

`ifndef __CACHE_TU_SVH__
`define __CACHE_TU_SVH__

typedef struct packed {
    logic __reserved;
} tu_op_req_t;

typedef struct packed {
    logic __reserved;
} tu_op_resp_t;

`endif

`endif