module hazard (
    ports
);
    
endmodule