//  Package: fetch_pkg
//
package fetch_pkg;
    import common::*;
    //  Group: Parameters
    

    //  Group: Typedefs
    typedef struct packed {
        word_t instr_;
        word_t pcplus8;
    } fetch_data_t;

    
endpackage: fetch_pkg
