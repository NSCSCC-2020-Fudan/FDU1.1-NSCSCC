// `include "mips.svh"
`include "instr_bus.svh"
`include "data_bus.svh"


// axi
module mycpu_top(
    input logic[5:0] ext_int,  //high active

    input logic aclk,
    input logic aresetn,   //low active

    output logic [3:0] arid,
    output logic [31:0] araddr,
    output logic [3:0] arlen,
    output logic [2 :0] arsize ,
    output logic [1 :0] arburst,
    output logic [1 :0] arlock ,
    output logic [3 :0] arcache,
    output logic [2 :0] arprot ,
    output logic        arvalid,
    input logic        arready,
    input logic [3 :0] rid    ,
    input logic [31:0] rdata  ,
    input logic [1 :0] rresp  ,
    input logic        rlast  ,
    input logic        rvalid ,
    output logic        rready ,
    output logic [3 :0] awid   ,
    output logic [31:0] awaddr ,
    output logic [3 :0] awlen  ,
    output logic [2 :0] awsize ,
    output logic [1 :0] awburst,
    output logic [1 :0] awlock ,
    output logic [3 :0] awcache,
    output logic [2 :0] awprot ,
    output logic        awvalid,
    input logic        awready,
    output logic [3 :0] wid    ,
    output logic [31:0] wdata  ,
    output logic [3 :0] wstrb  ,
    output logic        wlast  ,
    output logic        wvalid ,
    input logic        wready ,
    input logic [3 :0] bid    ,
    input logic [1 :0] bresp  ,
    input logic        bvalid ,
    output logic        bready ,

    //debug interface
    output logic[31:0] debug_wb_pc,
    output logic[3:0] debug_wb_rf_wen,
    output creg_addr_t debug_wb_rf_wnum,
    output word_t debug_wb_rf_wdata
);
    (*mark_debug = "true"*) ibus_req_t  icache_req;
    (*mark_debug = "true"*) ibus_resp_t icache_resp;
    (*mark_debug = "true"*) dbus_req_t  dcache_req,     uncached_req;
    (*mark_debug = "true"*) dbus_resp_t dcache_resp,    uncached_resp;
    (*mark_debug = "true"*) addr_t      imem_req_vaddr, dmem_req_vaddr;

    mycpu #(.DO_ADDR_TRANSLATION(0)) mycpu(
        .clk(aclk), .resetn(aresetn), .*
    );

    CacheLayer layer_inst(.*);
endmodule
