module interrupt(
);

endmodule