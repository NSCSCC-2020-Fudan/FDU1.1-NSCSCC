module bru 
    import common::*;
    import decode_pkg::*;(
    input word_t src1, src2,
    input decoded_op_t op,
    output logic branch_taken
);
    assign branch_taken = ;
endmodule