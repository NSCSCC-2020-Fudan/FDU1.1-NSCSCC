`ifndef __SBUFFER_SVH
`define __SBUFFER_SVH

`include "mips.svh"

`define SBUFFER_SIZE        'd8
`define SBUFFER_WIDTH       'd3

`endif
