`include "MIPS.h"

module BiMux(input logic [31: 0]
    );

endmodule