`ifndef __AXI3_COMMON_SVH
`define __AXI3_COMMON_SVH

typedef logic [3:0] nibble_t;
typedef logic [31:0] word_t;

`endif