//  Package: exc_pkg
//
package exc_pkg;
    //  Group: Parameters
    

    //  Group: Typedefs
    typedef enum logic[4:0] { NONE, INTERUPT, INSTR, LOAD, SAVE, BP, SYS } exception_info_t;

    
endpackage: exc_pkg
