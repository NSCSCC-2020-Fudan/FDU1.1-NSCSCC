//  Package: issue_pkg
//
package issue_pkg;
    import common::*;
    //  Group: Parameters


    //  Group: Typedefs

    
endpackage: issue_pkg
