//  Package: renaming_pkg
//
package renaming_pkg;
    //  Group: Parameters
    

    //  Group: Typedefs
    

    
endpackage: renaming_pkg
