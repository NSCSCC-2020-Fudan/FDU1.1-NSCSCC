`include "MIPS.svh"

module Hazard(
        input logic [4: 0] 
        output logic 
    );
endmodule