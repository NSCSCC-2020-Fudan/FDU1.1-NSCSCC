module free_list (
    
);
    import common::*;
    import free_list_pkg::*;

    // free list
    free_list_t list;
    
    // read

    // write
endmodule