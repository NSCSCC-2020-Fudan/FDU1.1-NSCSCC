`include "../interface.svh"
module datapath 
    import common::*;(
    
);
    
endmodule