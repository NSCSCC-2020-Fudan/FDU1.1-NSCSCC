`ifndef __EXECUTE_SVH
`define __EXECUTE_SVH

`include "global.svh"

typedef struct packed {
    
} exec_data_t;

`endif
