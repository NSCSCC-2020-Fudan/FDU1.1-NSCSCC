module ALUCL (
        input word_t a,
        output word_t b
    );
    always_comb begin
        priority case (1'b1)
            a[31]: b = 32'd0;
            a[30]: b = 32'd1;
            a[29]: b = 32'd2;
            a[28]: b = 32'd3;
            a[27]: b = 32'd4;
            a[26]: b = 32'd5;
            a[25]: b = 32'd6;
            a[24]: b = 32'd7;
            a[23]: b = 32'd8;
            a[22]: b = 32'd9;
            a[21]: b = 32'd10;
            a[20]: b = 32'd11;
            a[19]: b = 32'd12;
            a[18]: b = 32'd13;
            a[17]: b = 32'd14;
            a[16]: b = 32'd15;
            a[15]: b = 32'd16;
            a[14]: b = 32'd17;
            a[13]: b = 32'd18;
            a[12]: b = 32'd19;
            a[11]: b = 32'd20;
            a[10]: b = 32'd21;
            a[9]: b = 32'd22;
            a[8]: b = 32'd23;
            a[7]: b = 32'd24;
            a[6]: b = 32'd25;
            a[5]: b = 32'd26;
            a[4]: b = 32'd27;
            a[3]: b = 32'd28;
            a[2]: b = 32'd29;
            a[1]: b = 32'd30;
            a[0]: b = 32'd31;
            default : b = 32'd32;
        endcase
    end
endmodule