`define CACHE_WITHOUT_MIPS