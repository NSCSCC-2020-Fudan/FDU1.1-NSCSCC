`include "MIPS.h"

module Memory(
    
    );
endmodule
