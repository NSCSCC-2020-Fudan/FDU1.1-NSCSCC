`ifndef __CACHE_COMMON_SVH__
`define __CACHE_COMMON_SVH__

`include "defs.svh"
`include "axi.svh"
`include "cache_bus.svh"

`endif