// renaming aliasing table
module rat (
    
);
    import common::*;
    import rat_pkg::*;
    // table
    table_t mapping_table;

    // write

    // read
    
endmodule