`ifndef __INTERFACE_SVH
`define __INTERFACE_SVH



`endif
