module exception(
);

endmodule