`ifndef __AXI3_COMMON_SVH
`define __AXI3_COMMON_SVH

// nibble：半个字节
typedef logic [3:0] nibble_t;
typedef logic [31:0] word_t;

`endif