`ifndef __GLOBAL_SVH
`define __GLOBAL_SVH

typedef logic[31:0] word_t;
typedef logic[4:0] creg_addr_t;
typedef logic[16:0] halfword_t;

`define ZERO_EXT 1'b1
`define SIGN_EXT 1'b0
`endif
