// NOTE: set as "global include"

`ifndef DISABLE_DEFAULT_TU
`define DISABLE_DEFAULT_TU
`endif