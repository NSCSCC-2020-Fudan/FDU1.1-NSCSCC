`ifndef __MIPS_SVH
`define __MIPS_SVH

`include "global.svh"
`include "cp0.svh"
`include "exception.svh"
`include "decode.svh"
`include "execute.svh"
`include "fetch.svh"
`include "pcsource.svh"
`include "hazard.svh"
`include "memory.svh"
`include "hilo.svh"
`include "pipregs.svh"
`include "regfile.svh"
`include "writeback.svh"
`include "interface.svh"

`endif