`include "mips.svh"

module Decode (
    Dreg.out in,
    Ereg.in out,
    rfi.decode rf
);
    
endmodule

module MainDec (
    
);
    
endmodule

module ALUDec (
    
);
    
endmodule