module fetch (
    
);
    
endmodule