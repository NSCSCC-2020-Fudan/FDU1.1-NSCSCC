// address generate unit
module agu 
    import common::*;
    (
    
);
    vaddr_t addr;
    word_t data;
    
endmodule