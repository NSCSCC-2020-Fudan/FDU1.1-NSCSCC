module execute (
    Ereg_intf.out in,
    
);
    
endmodule