//  Package: exc_pkg
//
package exception_pkg;
    //  Group: Parameters
    

    //  Group: Typedefs
    typedef struct packed {
        logic interrupt;
        logic ri;
        logic instr;
        logic load;
        logic save;
        logic bp;
        logic sys;
    } exception_info_t;
    
endpackage: exception_pkg
