module commit 
    import common::*;
    import commit_pkg::*;(
    
);
    execute_data_t dataE;
    commit_data_t dataC;

    
endmodule