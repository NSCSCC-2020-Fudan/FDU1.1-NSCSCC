`include "mips.svh"

