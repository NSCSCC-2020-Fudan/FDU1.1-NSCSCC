`ifndef __MIPS_SVH
`define __MIPS_SVH



`endif

