`include "mips.svh"

module bpbdecode(
		word_t pc, instr,
		output word_t destpc
    );
    
endmodule
