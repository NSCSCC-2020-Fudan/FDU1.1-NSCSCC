//  Package: issue_pkg
//
package issue_pkg;
    //  Group: Parameters
    parameter ISSUE_WIDTH = 6; // maximum issue
    parameter MACHINE_WIDTH = 2; // maximum decode&renaming

    //  Group: Typedefs
    

    
endpackage: issue_pkg
