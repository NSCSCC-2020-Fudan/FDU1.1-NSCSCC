`include "MIPS.svh"

module exception(

    output Exception exception
);

endmodule