`ifndef __MEMORY_SVH
`define __MEMORY_SVH

typedef struct packed {
    
} mem_data_t;

`endif
