`ifndef __HAZARD_SVH
`define __HAZARD_SVH



`endif
