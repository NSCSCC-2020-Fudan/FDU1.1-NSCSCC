`include "shared.svh"

