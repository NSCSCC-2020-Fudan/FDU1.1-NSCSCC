module arf (
    
);
    logic word_t[AREG_NUM-1:0] regfile;
    
endmodule