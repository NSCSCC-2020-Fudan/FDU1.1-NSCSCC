module renaming (
    
);
    
endmodule