`ifndef __MEMORY_SVH
`define __MEMORY_SVH

interface RAM(output m_r_t read, output m_w_t write);
    
    modport in(output );
    modport out(input );
endinterface

`endif
