module memory (
    ports
);
    
endmodule