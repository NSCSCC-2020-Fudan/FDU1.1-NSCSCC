//  Package: decode_pkg
//
package decode_pkg;
    //  Group: Parameters
    

    //  Group: Typedefs
    

    
endpackage: decode_pkg
