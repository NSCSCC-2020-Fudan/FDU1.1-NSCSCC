//  Package: issue_pkg
//
package issue_pkg;
    import common::*;
    //  Group: Parameters


    //  Group: Typedefs
    typedef struct packed {
        logic en;
    } struct_name;

    
endpackage: issue_pkg
