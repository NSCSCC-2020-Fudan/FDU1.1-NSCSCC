module execute 
    import common::*;(
    
);
    
endmodule