`include "MIPS.h"

module WriteBack(
        input logic [4: 0] Rt, Rd,
        input logic [2: 0] Type, 
        input logic [2: 0] Move,
        input logic [4: 0] Memory,
        inout logic [31: 0] Result,
    );

    
    
endmodule
