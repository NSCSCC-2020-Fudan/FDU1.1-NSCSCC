`ifndef __PIPREGS_SVH
`define __PIPREGS_SVH

`include "mips.svh"

`endif
