`include "mips.svh"
module execute_ (
    decode_ereg_exec.exec in,
    exec_mreg_memory.exec out,
    hazard_intf.exec hazard
);
    word_t srca, srcb, srcb0;
    wrmux wrmux0(.rt(in.dataD.decoded_instr.rt), .rd(in.dataD.decoded_instr.rd), .jump(in.dataD.decoded_instr.ctl.jump), .regdst(in.dataD.decoded_instr.ctl.regdst), .writereg(out.dataE_new.writereg));
    srcaemux srcaemux(.e(in.dataD.srca),.m(hazard.aluoutM),.w(hazard.resultW),.sel(hazard.forwardAE),.srca);
    wdmux wdmux(.e(in.dataD.srcb),.m(hazard.aluoutM),.w(hazard.resultW),.sel(hazard.forwardBE),.srcb0);
    srcbemux srcbemux(.srcb0,.imm(in.dataD.decoded_instr.extended_imm),.shamt(in.dataD.decoded_instr.shamt),.srcb);
    alu alu(srca, srcb, in.dataD.decoded_instr.ctl.alufunc, out.dataE_new.aluout, out.dataE_new.exception_of);
    mult multdiv(.a(srca), .b(srcb), .op(in.dataD.decoded_instr.op), .hi(out.dataE_new.hi), .lo(out.dataE_new.lo));

    assign out.dataE_new.decoded_instr = in.dataD.decoded_instr;
    assign out.dataE_new.exception_instr = in.dataD.exception_instr;
    assign out.dataE_new.exception_ri = in.dataD.exception_ri;
    assign out.dataE_new.pcplus4 = in.dataD.pcplus4;
    assign hazard.dataE = out.dataE_new;
endmodule