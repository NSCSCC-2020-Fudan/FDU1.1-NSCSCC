`ifndef __WRITEDATA_SVH
`define __WRITEDATA_SVH

`define SB_W 8
`define SH_W 16

`endif
