//  Package: regfile_pkg
//
package regfile_pkg;
    //  Group: Parameters

    //  Group: Typedefs
    

    
endpackage: regfile_pkg
