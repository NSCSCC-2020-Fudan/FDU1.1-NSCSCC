`ifndef __MIPS_SVH
`define __MIPS_SVH

`include "global.svh"
`include "cp0.svh"
`include "exception.svh"
`include "pipregs.svh"
`include "pcsource.svh"
`include "regfile.svh"
`include "control.svh"

`endif

