`include "MIPS.h"

module Fetch(
        input logic clk,
        input logic [31: 0] PC,
        input logic [31: 0] RegJump, PCBranch, PCJump,
        input logic JumpReg, Branch, Jump,
    );

    

endmodule