module bru 
    import common::*;(
    input word_t src1, src2,
    input decode_pkg_t::decoded_op_t op
);
    
endmodule