`ifndef __WRITEBACK_SVH
`define __WRITEBACK_SVH



`endif
