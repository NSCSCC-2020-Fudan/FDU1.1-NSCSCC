module decode 
    import common::*;
    import decode_pkg::*;(
    
);
    
endmodule