//  Package: fetch_pkg
//
package fetch_pkg;
    import common::*;
    //  Group: Parameters
    

    //  Group: Typedefs
    

    
endpackage: fetch_pkg
